#misc abbreviations
#single upper case letter are usually initials
A
AB
B
C
D
E
F
G
H
I
J
K
L
M
N
O
P
Q
R
S
T
U
V
VG
W
X
Y
Z
dvs
etc
from
iaf
jfr
kl
kr
mao
mfl
mm
osv
pga
tex
tom
vs
